//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Sun Apr 25 13:44:04 2021
// Version: v12.5 12.900.10.16
//////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

// OSC_C0
module OSC_C0(
    // Inputs
    XTL,
    // Outputs
    XTLOSC_O2F
);

//--------------------------------------------------------------------
// Input
//--------------------------------------------------------------------
input  XTL;
//--------------------------------------------------------------------
// Output
//--------------------------------------------------------------------
output XTLOSC_O2F;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire   XTL;
wire   XTLOSC_O2F_net_0;
wire   XTLOSC_O2F_net_1;
//--------------------------------------------------------------------
// Top level output port assignments
//--------------------------------------------------------------------
assign XTLOSC_O2F_net_1 = XTLOSC_O2F_net_0;
assign XTLOSC_O2F       = XTLOSC_O2F_net_1;
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------OSC_C0_OSC_C0_0_OSC   -   Actel:SgCore:OSC:2.0.101
OSC_C0_OSC_C0_0_OSC OSC_C0_0(
        // Inputs
        .XTL                ( XTL ),
        // Outputs
        .RCOSC_25_50MHZ_CCC (  ),
        .RCOSC_25_50MHZ_O2F (  ),
        .RCOSC_1MHZ_CCC     (  ),
        .RCOSC_1MHZ_O2F     (  ),
        .XTLOSC_CCC         (  ),
        .XTLOSC_O2F         ( XTLOSC_O2F_net_0 ) 
        );


endmodule
